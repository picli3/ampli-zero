.title KiCad schematic
.include "/home/maykol/Documentos/spice/2SA1943.lib"
.include "/home/maykol/Documentos/spice/2SC5200.mod"
.include "/home/maykol/Documentos/spice/2n5401.lib"
.include "/home/maykol/Documentos/spice/2n5551.lib"
.include "/home/maykol/Documentos/spice/transistores_2.lib"
.save all
.probe alli
**comienzo de las pruebas
*.op
.tran 1u 5m 0
.measure tran Vo_RMS RMS v(/FB) from=0 to=1m
.measure tran Io_RMS RMS i(R112) from=0 to=1m
.measure tran Io_RMS(R101) RMS i(R101) from=0 to=5m

.meas tran skew5 FIND v(/FB) AT =0.75m

.control
	run
	plot (v(net-_q10-E_)- v(/FB))*i(R105)
	plot v(/FB)* i(r112)
	plot i(r101)*i(r101)*100
.endc

.control
	run
	tran 1u 5m 0
	print tran Io_RMS RMS v(vdb) from=0 to=1m
.endc


**
**.control
**fourier 1k v(/FB)
**gnuplot Vo v(/FB) v(/v4i)
**+ xycontour
**+ title 'Voltaje de salida Vs Voltaje de entrada'
**+ xlabel 'Tiempo (S)'
**+ ylabel 'Voltaje (V)'
**.endc

**Fin de las pruebas
*.tran 1u 5m 0
R13 /VB2 /gndv 10k
Q3 /VB2 Net-_Q3-B_ +32 2N5401
R14 /VE2 Net-_Q3-B_ 1k
R12 /gndv GND 12k
Q2 /VC2 /VB2 /VE2 2N5401
R9 +32 /VE2 150
Q7 Net-_Q4-C_ Net-_Q7-B_ Net-_Q7-E_ 2N5401
R18 /VC2 Net-_Q7-E_ 100
R22 Net-_Q7-B_ GND 10k
V1 +32 GND DC 32 
C102 Net-_Q7-B_ /v4i 3.3u
V4 /v4i GND DC 0 SIN( 0 1 1k 0 0 0 2 ) AC 2 
V2 GND -32 DC 32 
R15 Net-_Q5-E_ -32 68
Q5 Net-_Q4-B_ Net-_Q4-B_ Net-_Q5-E_ 2N5551
C7 Net-_C7-Pad1_ /FB 100p
R19 Net-_Q8-B_ Net-_C7-Pad1_ 220
R23 Net-_Q8-B_ /FB 18k
Q8 Net-_Q4-B_ Net-_Q8-B_ Net-_Q8-E_ 2N5401
R11 /VC2 Net-_Q8-E_ 100
R20 Net-_C6-Pad1_ Net-_Q8-B_ 1k
C6 Net-_C6-Pad1_ GND 220u
R10 Net-_Q4-E_ -32 68
Q4 Net-_Q4-C_ Net-_Q4-B_ Net-_Q4-E_ 2N5551
C8 -32 GND 100n
C3 +32 /gndv 10u
R101 +32 Net-_Q102-E_ 100
R115 /vdt Net-_Q112-B_ 1.2k
Q112 /vdt Net-_Q112-B_ vdb 2N5551
Q102 /vdt /VB2 Net-_Q102-E_ 2N5401
C5 Net-_Q4-C_ vdb 300p
R116 Net-_Q112-B_ vdb 330
Q9 vdb Net-_Q4-C_ Net-_Q9-E_ 2N5551
R21 Net-_Q9-E_ -32 22
R112 /FB Net-_L102-Pad1_ 6.4
R106 /FB Net-_Q101-E_ 0.33
Q10 +32 Net-_J2-Pin_1_ Net-_Q10-E_ 2SC5200
R105 Net-_Q10-E_ /FB 0.33
Q103 +32 /vdt Net-_J2-Pin_1_ 2SD669
R104 Net-_J2-Pin_1_ /FB 33
R103 /FB Net-_J3-Pin_1_ 33
XQ101 -32 Net-_J3-Pin_1_ Net-_Q101-E_ 2SA1943
Q104 -32 vdb Net-_J3-Pin_1_ 2SB649
C103 GND Net-_C103-Pad2_ 240u
R110 Net-_C103-Pad2_ GND 15
R111 Net-_L102-Pad1_ Net-_C103-Pad2_ 15
L102 Net-_L102-Pad1_ Net-_C103-Pad2_ 1m
L101 Net-_C103-Pad2_ GND 43m
.end
